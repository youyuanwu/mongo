module mongo

fn test_mongo_db(){
	assert 1 == 1
}